// DDR3AXI4.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module DDR3AXI4 (
		output wire        afi_half_clk_clk,                      //      afi_half_clk.clk
		output wire        afi_reset_reset_n,                     //         afi_reset.reset_n
		input  wire [3:0]  axi_translator_s0_awid,                // axi_translator_s0.awid
		input  wire [29:0] axi_translator_s0_awaddr,              //                  .awaddr
		input  wire [7:0]  axi_translator_s0_awlen,               //                  .awlen
		input  wire [2:0]  axi_translator_s0_awsize,              //                  .awsize
		input  wire [1:0]  axi_translator_s0_awburst,             //                  .awburst
		input  wire [0:0]  axi_translator_s0_awlock,              //                  .awlock
		input  wire [3:0]  axi_translator_s0_awcache,             //                  .awcache
		input  wire [2:0]  axi_translator_s0_awprot,              //                  .awprot
		input  wire [3:0]  axi_translator_s0_awqos,               //                  .awqos
		input  wire        axi_translator_s0_awvalid,             //                  .awvalid
		output wire        axi_translator_s0_awready,             //                  .awready
		input  wire [63:0] axi_translator_s0_wdata,               //                  .wdata
		input  wire [7:0]  axi_translator_s0_wstrb,               //                  .wstrb
		input  wire        axi_translator_s0_wlast,               //                  .wlast
		input  wire        axi_translator_s0_wvalid,              //                  .wvalid
		output wire        axi_translator_s0_wready,              //                  .wready
		output wire [3:0]  axi_translator_s0_bid,                 //                  .bid
		output wire [1:0]  axi_translator_s0_bresp,               //                  .bresp
		output wire        axi_translator_s0_bvalid,              //                  .bvalid
		input  wire        axi_translator_s0_bready,              //                  .bready
		input  wire [3:0]  axi_translator_s0_arid,                //                  .arid
		input  wire [29:0] axi_translator_s0_araddr,              //                  .araddr
		input  wire [7:0]  axi_translator_s0_arlen,               //                  .arlen
		input  wire [2:0]  axi_translator_s0_arsize,              //                  .arsize
		input  wire [1:0]  axi_translator_s0_arburst,             //                  .arburst
		input  wire [0:0]  axi_translator_s0_arlock,              //                  .arlock
		input  wire [3:0]  axi_translator_s0_arcache,             //                  .arcache
		input  wire [2:0]  axi_translator_s0_arprot,              //                  .arprot
		input  wire [3:0]  axi_translator_s0_arqos,               //                  .arqos
		input  wire        axi_translator_s0_arvalid,             //                  .arvalid
		output wire        axi_translator_s0_arready,             //                  .arready
		output wire [3:0]  axi_translator_s0_rid,                 //                  .rid
		output wire [63:0] axi_translator_s0_rdata,               //                  .rdata
		output wire [1:0]  axi_translator_s0_rresp,               //                  .rresp
		output wire        axi_translator_s0_rlast,               //                  .rlast
		output wire        axi_translator_s0_rvalid,              //                  .rvalid
		input  wire        axi_translator_s0_rready,              //                  .rready
		input  wire        clk_clk,                               //               clk.clk
		output wire [13:0] mem_mem_a,                             //               mem.mem_a
		output wire [2:0]  mem_mem_ba,                            //                  .mem_ba
		output wire [0:0]  mem_mem_ck,                            //                  .mem_ck
		output wire [0:0]  mem_mem_ck_n,                          //                  .mem_ck_n
		output wire [0:0]  mem_mem_cke,                           //                  .mem_cke
		output wire [0:0]  mem_mem_cs_n,                          //                  .mem_cs_n
		output wire [7:0]  mem_mem_dm,                            //                  .mem_dm
		output wire [0:0]  mem_mem_ras_n,                         //                  .mem_ras_n
		output wire [0:0]  mem_mem_cas_n,                         //                  .mem_cas_n
		output wire [0:0]  mem_mem_we_n,                          //                  .mem_we_n
		output wire        mem_mem_reset_n,                       //                  .mem_reset_n
		inout  wire [63:0] mem_mem_dq,                            //                  .mem_dq
		inout  wire [7:0]  mem_mem_dqs,                           //                  .mem_dqs
		inout  wire [7:0]  mem_mem_dqs_n,                         //                  .mem_dqs_n
		output wire [0:0]  mem_mem_odt,                           //                  .mem_odt
		input  wire        oct_rdn,                               //               oct.rdn
		input  wire        oct_rup,                               //                  .rup
		output wire        pll_sharing_pll_mem_clk,               //       pll_sharing.pll_mem_clk
		output wire        pll_sharing_pll_write_clk,             //                  .pll_write_clk
		output wire        pll_sharing_pll_locked,                //                  .pll_locked
		output wire        pll_sharing_pll_write_clk_pre_phy_clk, //                  .pll_write_clk_pre_phy_clk
		output wire        pll_sharing_pll_addr_cmd_clk,          //                  .pll_addr_cmd_clk
		output wire        pll_sharing_pll_avl_clk,               //                  .pll_avl_clk
		output wire        pll_sharing_pll_config_clk,            //                  .pll_config_clk
		input  wire        reset_reset_n                          //             reset.reset_n
	);

	wire    [1:0] merlin_axi_translator_0_m0_awburst;                          // merlin_axi_translator_0:m0_awburst -> mm_interconnect_0:merlin_axi_translator_0_m0_awburst
	wire    [7:0] merlin_axi_translator_0_m0_arlen;                            // merlin_axi_translator_0:m0_arlen -> mm_interconnect_0:merlin_axi_translator_0_m0_arlen
	wire    [3:0] merlin_axi_translator_0_m0_arqos;                            // merlin_axi_translator_0:m0_arqos -> mm_interconnect_0:merlin_axi_translator_0_m0_arqos
	wire    [7:0] merlin_axi_translator_0_m0_wstrb;                            // merlin_axi_translator_0:m0_wstrb -> mm_interconnect_0:merlin_axi_translator_0_m0_wstrb
	wire          merlin_axi_translator_0_m0_wready;                           // mm_interconnect_0:merlin_axi_translator_0_m0_wready -> merlin_axi_translator_0:m0_wready
	wire    [3:0] merlin_axi_translator_0_m0_rid;                              // mm_interconnect_0:merlin_axi_translator_0_m0_rid -> merlin_axi_translator_0:m0_rid
	wire          merlin_axi_translator_0_m0_rready;                           // merlin_axi_translator_0:m0_rready -> mm_interconnect_0:merlin_axi_translator_0_m0_rready
	wire    [7:0] merlin_axi_translator_0_m0_awlen;                            // merlin_axi_translator_0:m0_awlen -> mm_interconnect_0:merlin_axi_translator_0_m0_awlen
	wire    [3:0] merlin_axi_translator_0_m0_awqos;                            // merlin_axi_translator_0:m0_awqos -> mm_interconnect_0:merlin_axi_translator_0_m0_awqos
	wire    [3:0] merlin_axi_translator_0_m0_arcache;                          // merlin_axi_translator_0:m0_arcache -> mm_interconnect_0:merlin_axi_translator_0_m0_arcache
	wire          merlin_axi_translator_0_m0_wvalid;                           // merlin_axi_translator_0:m0_wvalid -> mm_interconnect_0:merlin_axi_translator_0_m0_wvalid
	wire   [29:0] merlin_axi_translator_0_m0_araddr;                           // merlin_axi_translator_0:m0_araddr -> mm_interconnect_0:merlin_axi_translator_0_m0_araddr
	wire    [2:0] merlin_axi_translator_0_m0_arprot;                           // merlin_axi_translator_0:m0_arprot -> mm_interconnect_0:merlin_axi_translator_0_m0_arprot
	wire    [2:0] merlin_axi_translator_0_m0_awprot;                           // merlin_axi_translator_0:m0_awprot -> mm_interconnect_0:merlin_axi_translator_0_m0_awprot
	wire   [63:0] merlin_axi_translator_0_m0_wdata;                            // merlin_axi_translator_0:m0_wdata -> mm_interconnect_0:merlin_axi_translator_0_m0_wdata
	wire          merlin_axi_translator_0_m0_arvalid;                          // merlin_axi_translator_0:m0_arvalid -> mm_interconnect_0:merlin_axi_translator_0_m0_arvalid
	wire    [3:0] merlin_axi_translator_0_m0_awcache;                          // merlin_axi_translator_0:m0_awcache -> mm_interconnect_0:merlin_axi_translator_0_m0_awcache
	wire    [3:0] merlin_axi_translator_0_m0_arid;                             // merlin_axi_translator_0:m0_arid -> mm_interconnect_0:merlin_axi_translator_0_m0_arid
	wire    [0:0] merlin_axi_translator_0_m0_arlock;                           // merlin_axi_translator_0:m0_arlock -> mm_interconnect_0:merlin_axi_translator_0_m0_arlock
	wire    [0:0] merlin_axi_translator_0_m0_awlock;                           // merlin_axi_translator_0:m0_awlock -> mm_interconnect_0:merlin_axi_translator_0_m0_awlock
	wire   [29:0] merlin_axi_translator_0_m0_awaddr;                           // merlin_axi_translator_0:m0_awaddr -> mm_interconnect_0:merlin_axi_translator_0_m0_awaddr
	wire    [1:0] merlin_axi_translator_0_m0_bresp;                            // mm_interconnect_0:merlin_axi_translator_0_m0_bresp -> merlin_axi_translator_0:m0_bresp
	wire          merlin_axi_translator_0_m0_arready;                          // mm_interconnect_0:merlin_axi_translator_0_m0_arready -> merlin_axi_translator_0:m0_arready
	wire   [63:0] merlin_axi_translator_0_m0_rdata;                            // mm_interconnect_0:merlin_axi_translator_0_m0_rdata -> merlin_axi_translator_0:m0_rdata
	wire          merlin_axi_translator_0_m0_awready;                          // mm_interconnect_0:merlin_axi_translator_0_m0_awready -> merlin_axi_translator_0:m0_awready
	wire    [1:0] merlin_axi_translator_0_m0_arburst;                          // merlin_axi_translator_0:m0_arburst -> mm_interconnect_0:merlin_axi_translator_0_m0_arburst
	wire    [2:0] merlin_axi_translator_0_m0_arsize;                           // merlin_axi_translator_0:m0_arsize -> mm_interconnect_0:merlin_axi_translator_0_m0_arsize
	wire          merlin_axi_translator_0_m0_bready;                           // merlin_axi_translator_0:m0_bready -> mm_interconnect_0:merlin_axi_translator_0_m0_bready
	wire          merlin_axi_translator_0_m0_rlast;                            // mm_interconnect_0:merlin_axi_translator_0_m0_rlast -> merlin_axi_translator_0:m0_rlast
	wire          merlin_axi_translator_0_m0_wlast;                            // merlin_axi_translator_0:m0_wlast -> mm_interconnect_0:merlin_axi_translator_0_m0_wlast
	wire    [1:0] merlin_axi_translator_0_m0_rresp;                            // mm_interconnect_0:merlin_axi_translator_0_m0_rresp -> merlin_axi_translator_0:m0_rresp
	wire    [3:0] merlin_axi_translator_0_m0_awid;                             // merlin_axi_translator_0:m0_awid -> mm_interconnect_0:merlin_axi_translator_0_m0_awid
	wire    [3:0] merlin_axi_translator_0_m0_bid;                              // mm_interconnect_0:merlin_axi_translator_0_m0_bid -> merlin_axi_translator_0:m0_bid
	wire          merlin_axi_translator_0_m0_bvalid;                           // mm_interconnect_0:merlin_axi_translator_0_m0_bvalid -> merlin_axi_translator_0:m0_bvalid
	wire    [2:0] merlin_axi_translator_0_m0_awsize;                           // merlin_axi_translator_0:m0_awsize -> mm_interconnect_0:merlin_axi_translator_0_m0_awsize
	wire          merlin_axi_translator_0_m0_awvalid;                          // merlin_axi_translator_0:m0_awvalid -> mm_interconnect_0:merlin_axi_translator_0_m0_awvalid
	wire          merlin_axi_translator_0_m0_rvalid;                           // mm_interconnect_0:merlin_axi_translator_0_m0_rvalid -> merlin_axi_translator_0:m0_rvalid
	wire          mm_interconnect_0_mem_if_ddr3_emif_0_avl_beginbursttransfer; // mm_interconnect_0:mem_if_ddr3_emif_0_avl_beginbursttransfer -> mem_if_ddr3_emif_0:avl_burstbegin
	wire  [255:0] mm_interconnect_0_mem_if_ddr3_emif_0_avl_readdata;           // mem_if_ddr3_emif_0:avl_rdata -> mm_interconnect_0:mem_if_ddr3_emif_0_avl_readdata
	wire          mm_interconnect_0_mem_if_ddr3_emif_0_avl_waitrequest;        // mem_if_ddr3_emif_0:avl_ready -> mm_interconnect_0:mem_if_ddr3_emif_0_avl_waitrequest
	wire   [24:0] mm_interconnect_0_mem_if_ddr3_emif_0_avl_address;            // mm_interconnect_0:mem_if_ddr3_emif_0_avl_address -> mem_if_ddr3_emif_0:avl_addr
	wire          mm_interconnect_0_mem_if_ddr3_emif_0_avl_read;               // mm_interconnect_0:mem_if_ddr3_emif_0_avl_read -> mem_if_ddr3_emif_0:avl_read_req
	wire   [31:0] mm_interconnect_0_mem_if_ddr3_emif_0_avl_byteenable;         // mm_interconnect_0:mem_if_ddr3_emif_0_avl_byteenable -> mem_if_ddr3_emif_0:avl_be
	wire          mm_interconnect_0_mem_if_ddr3_emif_0_avl_readdatavalid;      // mem_if_ddr3_emif_0:avl_rdata_valid -> mm_interconnect_0:mem_if_ddr3_emif_0_avl_readdatavalid
	wire          mm_interconnect_0_mem_if_ddr3_emif_0_avl_write;              // mm_interconnect_0:mem_if_ddr3_emif_0_avl_write -> mem_if_ddr3_emif_0:avl_write_req
	wire  [255:0] mm_interconnect_0_mem_if_ddr3_emif_0_avl_writedata;          // mm_interconnect_0:mem_if_ddr3_emif_0_avl_writedata -> mem_if_ddr3_emif_0:avl_wdata
	wire    [3:0] mm_interconnect_0_mem_if_ddr3_emif_0_avl_burstcount;         // mm_interconnect_0:mem_if_ddr3_emif_0_avl_burstcount -> mem_if_ddr3_emif_0:avl_size
	wire          mem_if_ddr3_emif_0_afi_clk_clk;                              // mem_if_ddr3_emif_0:afi_clk -> [mm_interconnect_0:mem_if_ddr3_emif_0_afi_clk_clk, rst_controller_001:clk]
	wire          rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [merlin_axi_translator_0:aresetn, mm_interconnect_0:merlin_axi_translator_0_clk_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [mm_interconnect_0:mem_if_ddr3_emif_0_avl_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:mem_if_ddr3_emif_0_soft_reset_reset_bridge_in_reset_reset]

	DDR3AXI4_mem_if_ddr3_emif_0 mem_if_ddr3_emif_0 (
		.pll_ref_clk               (clk_clk),                                                     //      pll_ref_clk.clk
		.global_reset_n            (reset_reset_n),                                               //     global_reset.reset_n
		.soft_reset_n              (reset_reset_n),                                               //       soft_reset.reset_n
		.afi_clk                   (mem_if_ddr3_emif_0_afi_clk_clk),                              //          afi_clk.clk
		.afi_half_clk              (afi_half_clk_clk),                                            //     afi_half_clk.clk
		.afi_reset_n               (afi_reset_reset_n),                                           //        afi_reset.reset_n
		.afi_reset_export_n        (),                                                            // afi_reset_export.reset_n
		.mem_a                     (mem_mem_a),                                                   //           memory.mem_a
		.mem_ba                    (mem_mem_ba),                                                  //                 .mem_ba
		.mem_ck                    (mem_mem_ck),                                                  //                 .mem_ck
		.mem_ck_n                  (mem_mem_ck_n),                                                //                 .mem_ck_n
		.mem_cke                   (mem_mem_cke),                                                 //                 .mem_cke
		.mem_cs_n                  (mem_mem_cs_n),                                                //                 .mem_cs_n
		.mem_dm                    (mem_mem_dm),                                                  //                 .mem_dm
		.mem_ras_n                 (mem_mem_ras_n),                                               //                 .mem_ras_n
		.mem_cas_n                 (mem_mem_cas_n),                                               //                 .mem_cas_n
		.mem_we_n                  (mem_mem_we_n),                                                //                 .mem_we_n
		.mem_reset_n               (mem_mem_reset_n),                                             //                 .mem_reset_n
		.mem_dq                    (mem_mem_dq),                                                  //                 .mem_dq
		.mem_dqs                   (mem_mem_dqs),                                                 //                 .mem_dqs
		.mem_dqs_n                 (mem_mem_dqs_n),                                               //                 .mem_dqs_n
		.mem_odt                   (mem_mem_odt),                                                 //                 .mem_odt
		.avl_ready                 (mm_interconnect_0_mem_if_ddr3_emif_0_avl_waitrequest),        //              avl.waitrequest_n
		.avl_burstbegin            (mm_interconnect_0_mem_if_ddr3_emif_0_avl_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr                  (mm_interconnect_0_mem_if_ddr3_emif_0_avl_address),            //                 .address
		.avl_rdata_valid           (mm_interconnect_0_mem_if_ddr3_emif_0_avl_readdatavalid),      //                 .readdatavalid
		.avl_rdata                 (mm_interconnect_0_mem_if_ddr3_emif_0_avl_readdata),           //                 .readdata
		.avl_wdata                 (mm_interconnect_0_mem_if_ddr3_emif_0_avl_writedata),          //                 .writedata
		.avl_be                    (mm_interconnect_0_mem_if_ddr3_emif_0_avl_byteenable),         //                 .byteenable
		.avl_read_req              (mm_interconnect_0_mem_if_ddr3_emif_0_avl_read),               //                 .read
		.avl_write_req             (mm_interconnect_0_mem_if_ddr3_emif_0_avl_write),              //                 .write
		.avl_size                  (mm_interconnect_0_mem_if_ddr3_emif_0_avl_burstcount),         //                 .burstcount
		.local_init_done           (),                                                            //           status.local_init_done
		.local_cal_success         (),                                                            //                 .local_cal_success
		.local_cal_fail            (),                                                            //                 .local_cal_fail
		.oct_rdn                   (oct_rdn),                                                     //              oct.rdn
		.oct_rup                   (oct_rup),                                                     //                 .rup
		.pll_mem_clk               (pll_sharing_pll_mem_clk),                                     //      pll_sharing.pll_mem_clk
		.pll_write_clk             (pll_sharing_pll_write_clk),                                   //                 .pll_write_clk
		.pll_locked                (pll_sharing_pll_locked),                                      //                 .pll_locked
		.pll_write_clk_pre_phy_clk (pll_sharing_pll_write_clk_pre_phy_clk),                       //                 .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk          (pll_sharing_pll_addr_cmd_clk),                                //                 .pll_addr_cmd_clk
		.pll_avl_clk               (pll_sharing_pll_avl_clk),                                     //                 .pll_avl_clk
		.pll_config_clk            (pll_sharing_pll_config_clk)                                   //                 .pll_config_clk
	);

	altera_merlin_axi_translator #(
		.USE_S0_AWID                       (1),
		.USE_S0_AWREGION                   (0),
		.USE_M0_AWREGION                   (0),
		.USE_S0_AWLEN                      (1),
		.USE_S0_AWSIZE                     (1),
		.USE_S0_AWBURST                    (1),
		.USE_S0_AWLOCK                     (1),
		.USE_M0_AWLOCK                     (1),
		.USE_S0_AWCACHE                    (1),
		.USE_M0_AWCACHE                    (1),
		.USE_M0_AWPROT                     (1),
		.USE_S0_AWQOS                      (1),
		.USE_M0_AWQOS                      (1),
		.USE_S0_WSTRB                      (1),
		.USE_M0_WLAST                      (1),
		.USE_S0_BID                        (1),
		.USE_S0_BRESP                      (1),
		.USE_M0_BRESP                      (1),
		.USE_S0_ARID                       (1),
		.USE_S0_ARREGION                   (0),
		.USE_M0_ARREGION                   (0),
		.USE_S0_ARLEN                      (1),
		.USE_S0_ARSIZE                     (1),
		.USE_S0_ARBURST                    (1),
		.USE_S0_ARLOCK                     (1),
		.USE_M0_ARLOCK                     (1),
		.USE_M0_ARCACHE                    (1),
		.USE_M0_ARQOS                      (1),
		.USE_M0_ARPROT                     (1),
		.USE_S0_ARCACHE                    (1),
		.USE_S0_ARQOS                      (1),
		.USE_S0_RID                        (1),
		.USE_S0_RRESP                      (1),
		.USE_M0_RRESP                      (1),
		.USE_S0_RLAST                      (1),
		.M0_ID_WIDTH                       (4),
		.DATA_WIDTH                        (64),
		.S0_ID_WIDTH                       (4),
		.M0_ADDR_WIDTH                     (30),
		.S0_WRITE_ADDR_USER_WIDTH          (64),
		.S0_READ_ADDR_USER_WIDTH           (64),
		.M0_WRITE_ADDR_USER_WIDTH          (64),
		.M0_READ_ADDR_USER_WIDTH           (64),
		.S0_WRITE_DATA_USER_WIDTH          (64),
		.S0_WRITE_RESPONSE_DATA_USER_WIDTH (64),
		.S0_READ_DATA_USER_WIDTH           (64),
		.M0_WRITE_DATA_USER_WIDTH          (64),
		.M0_WRITE_RESPONSE_DATA_USER_WIDTH (64),
		.M0_READ_DATA_USER_WIDTH           (64),
		.S0_ADDR_WIDTH                     (30),
		.USE_S0_AWUSER                     (0),
		.USE_S0_ARUSER                     (0),
		.USE_S0_WUSER                      (0),
		.USE_S0_RUSER                      (0),
		.USE_S0_BUSER                      (0),
		.USE_M0_AWUSER                     (0),
		.USE_M0_ARUSER                     (0),
		.USE_M0_WUSER                      (0),
		.USE_M0_RUSER                      (0),
		.USE_M0_BUSER                      (0),
		.M0_AXI_VERSION                    ("AXI4"),
		.M0_BURST_LENGTH_WIDTH             (8),
		.S0_BURST_LENGTH_WIDTH             (8),
		.M0_LOCK_WIDTH                     (1),
		.S0_LOCK_WIDTH                     (1),
		.S0_AXI_VERSION                    ("AXI4")
	) merlin_axi_translator_0 (
		.aclk        (afi_half_clk_clk),                                                              //       clk.clk
		.aresetn     (~rst_controller_reset_out_reset),                                      // clk_reset.reset_n
		.m0_awid     (merlin_axi_translator_0_m0_awid),                                      //        m0.awid
		.m0_awaddr   (merlin_axi_translator_0_m0_awaddr),                                    //          .awaddr
		.m0_awlen    (merlin_axi_translator_0_m0_awlen),                                     //          .awlen
		.m0_awsize   (merlin_axi_translator_0_m0_awsize),                                    //          .awsize
		.m0_awburst  (merlin_axi_translator_0_m0_awburst),                                   //          .awburst
		.m0_awlock   (merlin_axi_translator_0_m0_awlock),                                    //          .awlock
		.m0_awcache  (merlin_axi_translator_0_m0_awcache),                                   //          .awcache
		.m0_awprot   (merlin_axi_translator_0_m0_awprot),                                    //          .awprot
		.m0_awqos    (merlin_axi_translator_0_m0_awqos),                                     //          .awqos
		.m0_awvalid  (merlin_axi_translator_0_m0_awvalid),                                   //          .awvalid
		.m0_awready  (merlin_axi_translator_0_m0_awready),                                   //          .awready
		.m0_wdata    (merlin_axi_translator_0_m0_wdata),                                     //          .wdata
		.m0_wstrb    (merlin_axi_translator_0_m0_wstrb),                                     //          .wstrb
		.m0_wlast    (merlin_axi_translator_0_m0_wlast),                                     //          .wlast
		.m0_wvalid   (merlin_axi_translator_0_m0_wvalid),                                    //          .wvalid
		.m0_wready   (merlin_axi_translator_0_m0_wready),                                    //          .wready
		.m0_bid      (merlin_axi_translator_0_m0_bid),                                       //          .bid
		.m0_bresp    (merlin_axi_translator_0_m0_bresp),                                     //          .bresp
		.m0_bvalid   (merlin_axi_translator_0_m0_bvalid),                                    //          .bvalid
		.m0_bready   (merlin_axi_translator_0_m0_bready),                                    //          .bready
		.m0_arid     (merlin_axi_translator_0_m0_arid),                                      //          .arid
		.m0_araddr   (merlin_axi_translator_0_m0_araddr),                                    //          .araddr
		.m0_arlen    (merlin_axi_translator_0_m0_arlen),                                     //          .arlen
		.m0_arsize   (merlin_axi_translator_0_m0_arsize),                                    //          .arsize
		.m0_arburst  (merlin_axi_translator_0_m0_arburst),                                   //          .arburst
		.m0_arlock   (merlin_axi_translator_0_m0_arlock),                                    //          .arlock
		.m0_arcache  (merlin_axi_translator_0_m0_arcache),                                   //          .arcache
		.m0_arprot   (merlin_axi_translator_0_m0_arprot),                                    //          .arprot
		.m0_arqos    (merlin_axi_translator_0_m0_arqos),                                     //          .arqos
		.m0_arvalid  (merlin_axi_translator_0_m0_arvalid),                                   //          .arvalid
		.m0_arready  (merlin_axi_translator_0_m0_arready),                                   //          .arready
		.m0_rid      (merlin_axi_translator_0_m0_rid),                                       //          .rid
		.m0_rdata    (merlin_axi_translator_0_m0_rdata),                                     //          .rdata
		.m0_rresp    (merlin_axi_translator_0_m0_rresp),                                     //          .rresp
		.m0_rlast    (merlin_axi_translator_0_m0_rlast),                                     //          .rlast
		.m0_rvalid   (merlin_axi_translator_0_m0_rvalid),                                    //          .rvalid
		.m0_rready   (merlin_axi_translator_0_m0_rready),                                    //          .rready
		.s0_awid     (axi_translator_s0_awid),                                               //        s0.awid
		.s0_awaddr   (axi_translator_s0_awaddr),                                             //          .awaddr
		.s0_awlen    (axi_translator_s0_awlen),                                              //          .awlen
		.s0_awsize   (axi_translator_s0_awsize),                                             //          .awsize
		.s0_awburst  (axi_translator_s0_awburst),                                            //          .awburst
		.s0_awlock   (axi_translator_s0_awlock),                                             //          .awlock
		.s0_awcache  (axi_translator_s0_awcache),                                            //          .awcache
		.s0_awprot   (axi_translator_s0_awprot),                                             //          .awprot
		.s0_awqos    (axi_translator_s0_awqos),                                              //          .awqos
		.s0_awvalid  (axi_translator_s0_awvalid),                                            //          .awvalid
		.s0_awready  (axi_translator_s0_awready),                                            //          .awready
		.s0_wdata    (axi_translator_s0_wdata),                                              //          .wdata
		.s0_wstrb    (axi_translator_s0_wstrb),                                              //          .wstrb
		.s0_wlast    (axi_translator_s0_wlast),                                              //          .wlast
		.s0_wvalid   (axi_translator_s0_wvalid),                                             //          .wvalid
		.s0_wready   (axi_translator_s0_wready),                                             //          .wready
		.s0_bid      (axi_translator_s0_bid),                                                //          .bid
		.s0_bresp    (axi_translator_s0_bresp),                                              //          .bresp
		.s0_bvalid   (axi_translator_s0_bvalid),                                             //          .bvalid
		.s0_bready   (axi_translator_s0_bready),                                             //          .bready
		.s0_arid     (axi_translator_s0_arid),                                               //          .arid
		.s0_araddr   (axi_translator_s0_araddr),                                             //          .araddr
		.s0_arlen    (axi_translator_s0_arlen),                                              //          .arlen
		.s0_arsize   (axi_translator_s0_arsize),                                             //          .arsize
		.s0_arburst  (axi_translator_s0_arburst),                                            //          .arburst
		.s0_arlock   (axi_translator_s0_arlock),                                             //          .arlock
		.s0_arcache  (axi_translator_s0_arcache),                                            //          .arcache
		.s0_arprot   (axi_translator_s0_arprot),                                             //          .arprot
		.s0_arqos    (axi_translator_s0_arqos),                                              //          .arqos
		.s0_arvalid  (axi_translator_s0_arvalid),                                            //          .arvalid
		.s0_arready  (axi_translator_s0_arready),                                            //          .arready
		.s0_rid      (axi_translator_s0_rid),                                                //          .rid
		.s0_rdata    (axi_translator_s0_rdata),                                              //          .rdata
		.s0_rresp    (axi_translator_s0_rresp),                                              //          .rresp
		.s0_rlast    (axi_translator_s0_rlast),                                              //          .rlast
		.s0_rvalid   (axi_translator_s0_rvalid),                                             //          .rvalid
		.s0_rready   (axi_translator_s0_rready),                                             //          .rready
		.m0_awuser   (),                                                                     // (terminated)
		.m0_awregion (),                                                                     // (terminated)
		.m0_wuser    (),                                                                     // (terminated)
		.m0_buser    (64'b0000000000000000000000000000000000000000000000000000000000000000), // (terminated)
		.m0_aruser   (),                                                                     // (terminated)
		.m0_arregion (),                                                                     // (terminated)
		.m0_ruser    (64'b0000000000000000000000000000000000000000000000000000000000000000), // (terminated)
		.s0_awuser   (64'b0000000000000000000000000000000000000000000000000000000000000000), // (terminated)
		.s0_awregion (4'b0000),                                                              // (terminated)
		.s0_wuser    (64'b0000000000000000000000000000000000000000000000000000000000000000), // (terminated)
		.s0_buser    (),                                                                     // (terminated)
		.s0_aruser   (64'b0000000000000000000000000000000000000000000000000000000000000000), // (terminated)
		.s0_arregion (4'b0000),                                                              // (terminated)
		.s0_ruser    (),                                                                     // (terminated)
		.s0_wid      (4'b0000),                                                              // (terminated)
		.m0_wid      ()                                                                      // (terminated)
	);

	DDR3AXI4_mm_interconnect_0 mm_interconnect_0 (
		.merlin_axi_translator_0_m0_awid                                     (merlin_axi_translator_0_m0_awid),                             //                                    merlin_axi_translator_0_m0.awid
		.merlin_axi_translator_0_m0_awaddr                                   (merlin_axi_translator_0_m0_awaddr),                           //                                                              .awaddr
		.merlin_axi_translator_0_m0_awlen                                    (merlin_axi_translator_0_m0_awlen),                            //                                                              .awlen
		.merlin_axi_translator_0_m0_awsize                                   (merlin_axi_translator_0_m0_awsize),                           //                                                              .awsize
		.merlin_axi_translator_0_m0_awburst                                  (merlin_axi_translator_0_m0_awburst),                          //                                                              .awburst
		.merlin_axi_translator_0_m0_awlock                                   (merlin_axi_translator_0_m0_awlock),                           //                                                              .awlock
		.merlin_axi_translator_0_m0_awcache                                  (merlin_axi_translator_0_m0_awcache),                          //                                                              .awcache
		.merlin_axi_translator_0_m0_awprot                                   (merlin_axi_translator_0_m0_awprot),                           //                                                              .awprot
		.merlin_axi_translator_0_m0_awqos                                    (merlin_axi_translator_0_m0_awqos),                            //                                                              .awqos
		.merlin_axi_translator_0_m0_awvalid                                  (merlin_axi_translator_0_m0_awvalid),                          //                                                              .awvalid
		.merlin_axi_translator_0_m0_awready                                  (merlin_axi_translator_0_m0_awready),                          //                                                              .awready
		.merlin_axi_translator_0_m0_wdata                                    (merlin_axi_translator_0_m0_wdata),                            //                                                              .wdata
		.merlin_axi_translator_0_m0_wstrb                                    (merlin_axi_translator_0_m0_wstrb),                            //                                                              .wstrb
		.merlin_axi_translator_0_m0_wlast                                    (merlin_axi_translator_0_m0_wlast),                            //                                                              .wlast
		.merlin_axi_translator_0_m0_wvalid                                   (merlin_axi_translator_0_m0_wvalid),                           //                                                              .wvalid
		.merlin_axi_translator_0_m0_wready                                   (merlin_axi_translator_0_m0_wready),                           //                                                              .wready
		.merlin_axi_translator_0_m0_bid                                      (merlin_axi_translator_0_m0_bid),                              //                                                              .bid
		.merlin_axi_translator_0_m0_bresp                                    (merlin_axi_translator_0_m0_bresp),                            //                                                              .bresp
		.merlin_axi_translator_0_m0_bvalid                                   (merlin_axi_translator_0_m0_bvalid),                           //                                                              .bvalid
		.merlin_axi_translator_0_m0_bready                                   (merlin_axi_translator_0_m0_bready),                           //                                                              .bready
		.merlin_axi_translator_0_m0_arid                                     (merlin_axi_translator_0_m0_arid),                             //                                                              .arid
		.merlin_axi_translator_0_m0_araddr                                   (merlin_axi_translator_0_m0_araddr),                           //                                                              .araddr
		.merlin_axi_translator_0_m0_arlen                                    (merlin_axi_translator_0_m0_arlen),                            //                                                              .arlen
		.merlin_axi_translator_0_m0_arsize                                   (merlin_axi_translator_0_m0_arsize),                           //                                                              .arsize
		.merlin_axi_translator_0_m0_arburst                                  (merlin_axi_translator_0_m0_arburst),                          //                                                              .arburst
		.merlin_axi_translator_0_m0_arlock                                   (merlin_axi_translator_0_m0_arlock),                           //                                                              .arlock
		.merlin_axi_translator_0_m0_arcache                                  (merlin_axi_translator_0_m0_arcache),                          //                                                              .arcache
		.merlin_axi_translator_0_m0_arprot                                   (merlin_axi_translator_0_m0_arprot),                           //                                                              .arprot
		.merlin_axi_translator_0_m0_arqos                                    (merlin_axi_translator_0_m0_arqos),                            //                                                              .arqos
		.merlin_axi_translator_0_m0_arvalid                                  (merlin_axi_translator_0_m0_arvalid),                          //                                                              .arvalid
		.merlin_axi_translator_0_m0_arready                                  (merlin_axi_translator_0_m0_arready),                          //                                                              .arready
		.merlin_axi_translator_0_m0_rid                                      (merlin_axi_translator_0_m0_rid),                              //                                                              .rid
		.merlin_axi_translator_0_m0_rdata                                    (merlin_axi_translator_0_m0_rdata),                            //                                                              .rdata
		.merlin_axi_translator_0_m0_rresp                                    (merlin_axi_translator_0_m0_rresp),                            //                                                              .rresp
		.merlin_axi_translator_0_m0_rlast                                    (merlin_axi_translator_0_m0_rlast),                            //                                                              .rlast
		.merlin_axi_translator_0_m0_rvalid                                   (merlin_axi_translator_0_m0_rvalid),                           //                                                              .rvalid
		.merlin_axi_translator_0_m0_rready                                   (merlin_axi_translator_0_m0_rready),                           //                                                              .rready
		.clk_0_clk_clk                                                       (afi_half_clk_clk),                                                     //                                                     clk_0_clk.clk
		.mem_if_ddr3_emif_0_afi_clk_clk                                      (mem_if_ddr3_emif_0_afi_clk_clk),                              //                                    mem_if_ddr3_emif_0_afi_clk.clk
		.mem_if_ddr3_emif_0_avl_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // mem_if_ddr3_emif_0_avl_translator_reset_reset_bridge_in_reset.reset
		.mem_if_ddr3_emif_0_soft_reset_reset_bridge_in_reset_reset           (rst_controller_001_reset_out_reset),                          //           mem_if_ddr3_emif_0_soft_reset_reset_bridge_in_reset.reset
		.merlin_axi_translator_0_clk_reset_reset_bridge_in_reset_reset       (rst_controller_reset_out_reset),                              //       merlin_axi_translator_0_clk_reset_reset_bridge_in_reset.reset
		.mem_if_ddr3_emif_0_avl_address                                      (mm_interconnect_0_mem_if_ddr3_emif_0_avl_address),            //                                        mem_if_ddr3_emif_0_avl.address
		.mem_if_ddr3_emif_0_avl_write                                        (mm_interconnect_0_mem_if_ddr3_emif_0_avl_write),              //                                                              .write
		.mem_if_ddr3_emif_0_avl_read                                         (mm_interconnect_0_mem_if_ddr3_emif_0_avl_read),               //                                                              .read
		.mem_if_ddr3_emif_0_avl_readdata                                     (mm_interconnect_0_mem_if_ddr3_emif_0_avl_readdata),           //                                                              .readdata
		.mem_if_ddr3_emif_0_avl_writedata                                    (mm_interconnect_0_mem_if_ddr3_emif_0_avl_writedata),          //                                                              .writedata
		.mem_if_ddr3_emif_0_avl_beginbursttransfer                           (mm_interconnect_0_mem_if_ddr3_emif_0_avl_beginbursttransfer), //                                                              .beginbursttransfer
		.mem_if_ddr3_emif_0_avl_burstcount                                   (mm_interconnect_0_mem_if_ddr3_emif_0_avl_burstcount),         //                                                              .burstcount
		.mem_if_ddr3_emif_0_avl_byteenable                                   (mm_interconnect_0_mem_if_ddr3_emif_0_avl_byteenable),         //                                                              .byteenable
		.mem_if_ddr3_emif_0_avl_readdatavalid                                (mm_interconnect_0_mem_if_ddr3_emif_0_avl_readdatavalid),      //                                                              .readdatavalid
		.mem_if_ddr3_emif_0_avl_waitrequest                                  (~mm_interconnect_0_mem_if_ddr3_emif_0_avl_waitrequest)        //                                                              .waitrequest
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (mem_if_ddr3_emif_0_afi_clk_clk),     //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
